/*

Copyright (c) 2014-2021 Alex Forencich

Permission is hereby granted, free of charge, to any person obtaining a copy
of this software and associated documentation files (the "Software"), to deal
in the Software without restriction, including without limitation the rights
to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
copies of the Software, and to permit persons to whom the Software is
furnished to do so, subject to the following conditions:

The above copyright notice and this permission notice shall be included in
all copies or substantial portions of the Software.

THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY
FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
THE SOFTWARE.

*/

// Language: Verilog 2001

`include "config.vh"

`resetall
`default_nettype none

/*
 * AXI4-Stream asynchronous FIFO
 */
module axis_async_fifo #
(
    // FIFO depth in words
    // KEEP_WIDTH words per cycle if KEEP_ENABLE set
    // Rounded up to nearest power of 2 cycles
    parameter DEPTH = 4096,
    // Width of AXI stream interfaces in bits
    parameter DATA_WIDTH = 8,
    // Propagate tkeep signal
    // If disabled, tkeep assumed to be 1'b1
    parameter KEEP_ENABLE = (DATA_WIDTH>8),
    // tkeep signal width (words per cycle)
    parameter KEEP_WIDTH = ((DATA_WIDTH+7)/8),
    // Propagate tlast signal
    parameter LAST_ENABLE = 1,
    // Propagate tid signal
    parameter ID_ENABLE = 0,
    // tid signal width
    parameter ID_WIDTH = 8,
    // Propagate tdest signal
    parameter DEST_ENABLE = 0,
    // tdest signal width
    parameter DEST_WIDTH = 8,
    // Propagate tuser signal
    parameter USER_ENABLE = 1,
    // tuser signal width
    parameter USER_WIDTH = 1,
    // number of output pipeline registers
    parameter PIPELINE_OUTPUT = 2,
    // Frame FIFO mode - operate on frames instead of cycles
    // When set, m_axis_tvalid will not be deasserted within a frame
    // Requires LAST_ENABLE set
    parameter FRAME_FIFO = 0,
    // tuser value for bad frame marker
    parameter USER_BAD_FRAME_VALUE = 1'b1,
    // tuser mask for bad frame marker
    parameter USER_BAD_FRAME_MASK = 1'b1,
    // Drop frames larger than FIFO
    // Requires FRAME_FIFO set
    parameter DROP_OVERSIZE_FRAME = FRAME_FIFO,
    // Drop frames marked bad
    // Requires FRAME_FIFO and DROP_OVERSIZE_FRAME set
    parameter DROP_BAD_FRAME = 0,
    // Drop incoming frames when full
    // When set, s_axis_tready is always asserted
    // Requires FRAME_FIFO and DROP_OVERSIZE_FRAME set
    parameter DROP_WHEN_FULL = 0
)
(
    /*
     * AXI input
     */
    input  wire                   s_clk,
    input  wire                   s_rst_n,
    input  wire                   s_drop,
    input  wire [DATA_WIDTH-1:0]  s_axis_tdata,
    input  wire [KEEP_WIDTH-1:0]  s_axis_tkeep,
    input  wire                   s_axis_tvalid,
    output wire                   s_axis_tready,
    input  wire                   s_axis_tlast,
    input  wire [ID_WIDTH-1:0]    s_axis_tid,
    input  wire [DEST_WIDTH-1:0]  s_axis_tdest,
    input  wire [USER_WIDTH-1:0]  s_axis_tuser,

    /*
     * AXI output
     */
    input  wire                   m_clk,
    input  wire                   m_rst_n,
    output wire [DATA_WIDTH-1:0]  m_axis_tdata,
    output wire [KEEP_WIDTH-1:0]  m_axis_tkeep,
    output wire                   m_axis_tvalid,
    input  wire                   m_axis_tready,
    output wire                   m_axis_tlast,
    output wire [ID_WIDTH-1:0]    m_axis_tid,
    output wire [DEST_WIDTH-1:0]  m_axis_tdest,
    output wire [USER_WIDTH-1:0]  m_axis_tuser,

    /*
     * Status
     */
    output wire                   s_status_overflow,
    output wire                   s_status_bad_frame,
    output wire                   s_status_good_frame,
    output wire                   m_status_overflow,
    output wire                   m_status_bad_frame,
    output wire                   m_status_good_frame
);

localparam ADDR_WIDTH = (KEEP_ENABLE && KEEP_WIDTH > 1) ? $clog2(DEPTH/KEEP_WIDTH) : $clog2(DEPTH);

// check configuration
`ifdef TARGET_SIM
initial begin
    if (PIPELINE_OUTPUT < 1) begin
        $error("Error: PIPELINE_OUTPUT must be at least 1 (instance %m)");
        $finish;
    end

    if (FRAME_FIFO && !LAST_ENABLE) begin
        $error("Error: FRAME_FIFO set requires LAST_ENABLE set (instance %m)");
        $finish;
    end

    if (DROP_OVERSIZE_FRAME && !FRAME_FIFO) begin
        $error("Error: DROP_OVERSIZE_FRAME set requires FRAME_FIFO set (instance %m)");
        $finish;
    end

    if (DROP_BAD_FRAME && !(FRAME_FIFO && DROP_OVERSIZE_FRAME)) begin
        $error("Error: DROP_BAD_FRAME set requires FRAME_FIFO and DROP_OVERSIZE_FRAME set (instance %m)");
        $finish;
    end

    if (DROP_WHEN_FULL && !(FRAME_FIFO && DROP_OVERSIZE_FRAME)) begin
        $error("Error: DROP_WHEN_FULL set requires FRAME_FIFO and DROP_OVERSIZE_FRAME set (instance %m)");
        $finish;
    end

    if (DROP_BAD_FRAME && (USER_BAD_FRAME_MASK & {USER_WIDTH{1'b1}}) == 0) begin
        $error("Error: Invalid USER_BAD_FRAME_MASK value (instance %m)");
        $finish;
    end
end
`endif

localparam KEEP_OFFSET = DATA_WIDTH;
localparam LAST_OFFSET = KEEP_OFFSET + (KEEP_ENABLE ? KEEP_WIDTH : 0);
localparam ID_OFFSET   = LAST_OFFSET + (LAST_ENABLE ? 1          : 0);
localparam DEST_OFFSET = ID_OFFSET   + (ID_ENABLE   ? ID_WIDTH   : 0);
localparam USER_OFFSET = DEST_OFFSET + (DEST_ENABLE ? DEST_WIDTH : 0);
localparam WIDTH       = USER_OFFSET + (USER_ENABLE ? USER_WIDTH : 0);

reg [ADDR_WIDTH:0] wr_ptr_reg;
reg [ADDR_WIDTH:0] wr_ptr_cur_reg;
reg [ADDR_WIDTH:0] wr_ptr_gray_reg;
reg [ADDR_WIDTH:0] wr_ptr_sync_gray_reg;
reg [ADDR_WIDTH:0] wr_ptr_cur_gray_reg;
reg [ADDR_WIDTH:0] rd_ptr_reg;
reg [ADDR_WIDTH:0] rd_ptr_gray_reg;

(* SHREG_EXTRACT = "NO" *)
reg [ADDR_WIDTH:0] wr_ptr_gray_sync1_reg;
(* SHREG_EXTRACT = "NO" *)
reg [ADDR_WIDTH:0] wr_ptr_gray_sync2_reg;
(* SHREG_EXTRACT = "NO" *)
reg [ADDR_WIDTH:0] rd_ptr_gray_sync1_reg;
(* SHREG_EXTRACT = "NO" *)
reg [ADDR_WIDTH:0] rd_ptr_gray_sync2_reg;

reg wr_ptr_update_valid_reg;
reg wr_ptr_update_reg;
(* SHREG_EXTRACT = "NO" *)
reg wr_ptr_update_sync1_reg;
(* SHREG_EXTRACT = "NO" *)
reg wr_ptr_update_sync2_reg;
(* SHREG_EXTRACT = "NO" *)
reg wr_ptr_update_sync3_reg;
(* SHREG_EXTRACT = "NO" *)
reg wr_ptr_update_ack_sync1_reg;
(* SHREG_EXTRACT = "NO" *)
reg wr_ptr_update_ack_sync2_reg;

(* SHREG_EXTRACT = "NO" *)
reg s_rst_sync1_reg;
(* SHREG_EXTRACT = "NO" *)
reg s_rst_sync2_reg;
(* SHREG_EXTRACT = "NO" *)
reg s_rst_sync3_reg;
(* SHREG_EXTRACT = "NO" *)
reg m_rst_sync1_reg;
(* SHREG_EXTRACT = "NO" *)
reg m_rst_sync2_reg;
(* SHREG_EXTRACT = "NO" *)
reg m_rst_sync3_reg;

(* ramstyle = "no_rw_check" *)
reg [WIDTH-1:0] mem[(2**ADDR_WIDTH)-1:0];

wire [WIDTH-1:0] s_axis;

reg [WIDTH-1:0] m_axis_pipe_reg[PIPELINE_OUTPUT-1:0];
reg [PIPELINE_OUTPUT-1:0] m_axis_tvalid_pipe_reg;

// full when first TWO MSBs do NOT match, but rest matches
// (gray code equivalent of first MSB different but rest same)
wire full = wr_ptr_gray_reg == (rd_ptr_gray_sync2_reg ^ {2'b11, {ADDR_WIDTH-1{1'b0}}});
wire full_cur = wr_ptr_cur_gray_reg == (rd_ptr_gray_sync2_reg ^ {2'b11, {ADDR_WIDTH-1{1'b0}}});
// empty when pointers match exactly
wire empty = rd_ptr_gray_reg == (FRAME_FIFO ? wr_ptr_gray_sync1_reg : wr_ptr_gray_sync2_reg);
// overflow within packet
wire full_wr = wr_ptr_reg == (wr_ptr_cur_reg ^ {1'b1, {ADDR_WIDTH{1'b0}}});

reg s_frame_reg;
reg m_frame_reg;

reg drop_frame_reg;
reg send_frame_reg;
reg overflow_reg;
reg bad_frame_reg;
reg good_frame_reg;

reg m_drop_frame_reg;
reg m_terminate_frame_reg;

reg overflow_sync1_reg;
reg overflow_sync2_reg;
reg overflow_sync3_reg;
reg overflow_sync4_reg;
reg bad_frame_sync1_reg;
reg bad_frame_sync2_reg;
reg bad_frame_sync3_reg;
reg bad_frame_sync4_reg;
reg good_frame_sync1_reg;
reg good_frame_sync2_reg;
reg good_frame_sync3_reg;
reg good_frame_sync4_reg;

assign s_axis_tready = (FRAME_FIFO ? (!full_cur || (full_wr && DROP_OVERSIZE_FRAME) || DROP_WHEN_FULL) : !full) && s_rst_sync3_reg;

generate
    assign s_axis[DATA_WIDTH-1:0] = s_axis_tdata;
    if (KEEP_ENABLE) assign s_axis[KEEP_OFFSET +: KEEP_WIDTH] = s_axis_tkeep;
    if (LAST_ENABLE) assign s_axis[LAST_OFFSET]               = s_axis_tlast;
    if (ID_ENABLE)   assign s_axis[ID_OFFSET   +: ID_WIDTH]   = s_axis_tid;
    if (DEST_ENABLE) assign s_axis[DEST_OFFSET +: DEST_WIDTH] = s_axis_tdest;
    if (USER_ENABLE) assign s_axis[USER_OFFSET +: USER_WIDTH] = s_axis_tuser;
endgenerate

wire                   m_axis_tvalid_pipe = m_axis_tvalid_pipe_reg[PIPELINE_OUTPUT-1];

wire [DATA_WIDTH-1:0]  m_axis_tdata_pipe  = m_axis_pipe_reg[PIPELINE_OUTPUT-1][DATA_WIDTH-1:0];
wire [KEEP_WIDTH-1:0]  m_axis_tkeep_pipe  = KEEP_ENABLE ? m_axis_pipe_reg[PIPELINE_OUTPUT-1][KEEP_OFFSET +: KEEP_WIDTH] : {KEEP_WIDTH{1'b1}};
wire                   m_axis_tlast_pipe  = LAST_ENABLE ? m_axis_pipe_reg[PIPELINE_OUTPUT-1][LAST_OFFSET] : 1'b1;
wire [ID_WIDTH-1:0]    m_axis_tid_pipe    = ID_ENABLE   ? m_axis_pipe_reg[PIPELINE_OUTPUT-1][ID_OFFSET +: ID_WIDTH] : {ID_WIDTH{1'b0}};
wire [DEST_WIDTH-1:0]  m_axis_tdest_pipe  = DEST_ENABLE ? m_axis_pipe_reg[PIPELINE_OUTPUT-1][DEST_OFFSET +: DEST_WIDTH] : {DEST_WIDTH{1'b0}};
wire [USER_WIDTH-1:0]  m_axis_tuser_pipe  = USER_ENABLE ? m_axis_pipe_reg[PIPELINE_OUTPUT-1][USER_OFFSET +: USER_WIDTH] : {USER_WIDTH{1'b0}};

assign m_axis_tvalid = m_axis_tvalid_pipe;

assign m_axis_tdata = m_axis_tdata_pipe;
assign m_axis_tkeep = m_axis_tkeep_pipe;
assign m_axis_tlast = (m_terminate_frame_reg ? 1'b1 : m_axis_tlast_pipe);
assign m_axis_tid   = m_axis_tid_pipe;
assign m_axis_tdest = m_axis_tdest_pipe;
assign m_axis_tuser = (m_terminate_frame_reg ? USER_BAD_FRAME_VALUE : m_axis_tuser_pipe);

assign s_status_overflow = overflow_reg;
assign s_status_bad_frame = bad_frame_reg;
assign s_status_good_frame = good_frame_reg;

assign m_status_overflow = overflow_sync3_reg ^ overflow_sync4_reg;
assign m_status_bad_frame = bad_frame_sync3_reg ^ bad_frame_sync4_reg;
assign m_status_good_frame = good_frame_sync3_reg ^ good_frame_sync4_reg;

// reset synchronization
always @(posedge m_clk or negedge m_rst_n) begin
    if (!m_rst_n) begin
        s_rst_sync1_reg <= 1'b0;
    end else begin
        s_rst_sync1_reg <= 1'b1;
    end
end

always @(posedge s_clk or negedge s_rst_n) begin
    if (!s_rst_n) begin
        s_rst_sync2_reg <= 1'b0;
        s_rst_sync3_reg <= 1'b0;
    end else begin
        s_rst_sync2_reg <= s_rst_sync1_reg;
        s_rst_sync3_reg <= s_rst_sync2_reg;
    end
end

always @(posedge s_clk or negedge s_rst_n) begin
    if (!s_rst_n) begin
        m_rst_sync1_reg <= 1'b0;
    end else begin
        m_rst_sync1_reg <= 1'b1;
    end
end

always @(posedge m_clk or negedge m_rst_n) begin
    if (!m_rst_n) begin
        m_rst_sync2_reg <= 1'b0;
        m_rst_sync3_reg <= 1'b0;
    end else begin
        m_rst_sync2_reg <= m_rst_sync1_reg;
        m_rst_sync3_reg <= m_rst_sync2_reg;
    end
end

integer i;

// Write logic
`ifdef TARGET_XILINX
always @(posedge s_clk) begin // Vivado could not infer BRAM if async reset is used.
`else
always @(posedge s_clk or negedge s_rst_n) begin
`endif
    if (!s_rst_n) begin
`ifndef TARGET_XILINX
        for (i=0; i<(2**ADDR_WIDTH); i=i+1) begin
`ifdef TARGET_SIM
            mem[i] = 0;
`else
            mem[i] <= 0;
`endif
        end
`endif

        wr_ptr_reg <= {ADDR_WIDTH+1{1'b0}};
        wr_ptr_cur_reg <= {ADDR_WIDTH+1{1'b0}};
        wr_ptr_gray_reg <= {ADDR_WIDTH+1{1'b0}};
        wr_ptr_sync_gray_reg <= {ADDR_WIDTH+1{1'b0}};
        wr_ptr_cur_gray_reg <= {ADDR_WIDTH+1{1'b0}};

        wr_ptr_update_valid_reg <= 1'b0;
        wr_ptr_update_reg <= 1'b0;

        s_frame_reg <= 1'b0;

        drop_frame_reg <= 1'b0;
        send_frame_reg <= 1'b0;
        overflow_reg <= 1'b0;
        bad_frame_reg <= 1'b0;
        good_frame_reg <= 1'b0;
    end else begin
        overflow_reg <= 1'b0;
        bad_frame_reg <= 1'b0;
        good_frame_reg <= 1'b0;

        if (FRAME_FIFO && wr_ptr_update_valid_reg) begin
            // have updated pointer to sync
            if (wr_ptr_update_reg == wr_ptr_update_ack_sync2_reg) begin
                // no sync in progress; sync update
                wr_ptr_update_valid_reg <= 1'b0;
                wr_ptr_sync_gray_reg <= wr_ptr_gray_reg;
                wr_ptr_update_reg <= !wr_ptr_update_ack_sync2_reg;
            end
        end

        if (s_axis_tready && s_axis_tvalid && LAST_ENABLE) begin
            // track input frame status
            s_frame_reg <= !s_axis_tlast;
        end

        if (!s_rst_sync3_reg && LAST_ENABLE) begin
            // if sink side is reset during transfer, drop partial frame
            if (s_frame_reg && !(s_axis_tready && s_axis_tvalid && s_axis_tlast)) begin
                drop_frame_reg <= 1'b1;
            end
            if (s_axis_tready && s_axis_tvalid && !s_axis_tlast) begin
                drop_frame_reg <= 1'b1;
            end
        end

        if (s_axis_tready && s_axis_tvalid) begin
            // transfer in
            if (s_drop) begin
                drop_frame_reg <= 1;
            end
            if (!FRAME_FIFO) begin
                // normal FIFO mode
                mem[wr_ptr_reg[ADDR_WIDTH-1:0]] <= s_axis;
                if (drop_frame_reg && LAST_ENABLE) begin
                    // currently dropping frame
                    // (only for frame transfers interrupted by sink reset)
                    if (s_axis_tlast) begin
                        // end of frame, clear drop flag
                        drop_frame_reg <= s_drop;
                    end
                end else begin
                    // update pointers
                    wr_ptr_reg <= (wr_ptr_reg + 1);
                    wr_ptr_gray_reg <= (wr_ptr_reg + 1) ^ ((wr_ptr_reg + 1) >> 1);
                end
            end else if ((full_cur && DROP_WHEN_FULL) || (full_wr && DROP_OVERSIZE_FRAME) || drop_frame_reg) begin
                // full, packet overflow, or currently dropping frame
                // drop frame
                drop_frame_reg <= 1'b1;
                if (s_axis_tlast) begin
                    // end of frame, reset write pointer
                    wr_ptr_cur_reg <= wr_ptr_reg;
                    wr_ptr_cur_gray_reg <= wr_ptr_reg ^ (wr_ptr_reg >> 1);
                    drop_frame_reg <= s_drop;
                    overflow_reg <= 1'b1;
                end
            end else begin
                mem[wr_ptr_cur_reg[ADDR_WIDTH-1:0]] <= s_axis;
                wr_ptr_cur_reg <= wr_ptr_cur_reg + 1;
                wr_ptr_cur_gray_reg <= (wr_ptr_cur_reg + 1) ^ ((wr_ptr_cur_reg + 1) >> 1);
                if (s_axis_tlast || (!DROP_OVERSIZE_FRAME && (full_wr || send_frame_reg))) begin
                    // end of frame or send frame
                    send_frame_reg <= !s_axis_tlast;
                    if (s_axis_tlast && DROP_BAD_FRAME && USER_BAD_FRAME_MASK & ~(s_axis_tuser ^ USER_BAD_FRAME_VALUE)) begin
                        // bad packet, reset write pointer
                        wr_ptr_cur_reg <= wr_ptr_reg;
                        wr_ptr_cur_gray_reg <= wr_ptr_reg ^ (wr_ptr_reg >> 1);
                        bad_frame_reg <= 1'b1;
                    end else begin
                        // good packet or packet overflow, update write pointer
                        wr_ptr_reg <= wr_ptr_cur_reg + 1;
                        wr_ptr_gray_reg <= (wr_ptr_cur_reg + 1) ^ ((wr_ptr_cur_reg + 1) >> 1);

                        if (wr_ptr_update_reg == wr_ptr_update_ack_sync2_reg) begin
                            // no sync in progress; sync update
                            wr_ptr_update_valid_reg <= 1'b0;
                            wr_ptr_sync_gray_reg <= (wr_ptr_cur_reg + 1) ^ ((wr_ptr_cur_reg + 1) >> 1);
                            wr_ptr_update_reg <= !wr_ptr_update_ack_sync2_reg;
                        end else begin
                            // sync in progress; flag it for later
                            wr_ptr_update_valid_reg <= 1'b1;
                        end

                        good_frame_reg <= s_axis_tlast;
                    end
                end
            end
        end else if (s_axis_tvalid && full_wr && FRAME_FIFO && !DROP_OVERSIZE_FRAME) begin
            // data valid with packet overflow
            // update write pointer
            send_frame_reg <= 1'b1;
            wr_ptr_reg <= wr_ptr_cur_reg;
            wr_ptr_gray_reg <= wr_ptr_cur_reg ^ (wr_ptr_cur_reg >> 1);

            if (wr_ptr_update_reg == wr_ptr_update_ack_sync2_reg) begin
                // no sync in progress; sync update
                wr_ptr_update_valid_reg <= 1'b0;
                wr_ptr_sync_gray_reg <= wr_ptr_cur_reg ^ (wr_ptr_cur_reg >> 1);
                wr_ptr_update_reg <= !wr_ptr_update_ack_sync2_reg;
            end else begin
                // sync in progress; flag it for later
                wr_ptr_update_valid_reg <= 1'b1;
            end
        end

        if (!s_rst_sync3_reg) begin
            wr_ptr_reg <= {ADDR_WIDTH+1{1'b0}};
            wr_ptr_cur_reg <= {ADDR_WIDTH+1{1'b0}};
            wr_ptr_gray_reg <= {ADDR_WIDTH+1{1'b0}};
            wr_ptr_sync_gray_reg <= {ADDR_WIDTH+1{1'b0}};
            wr_ptr_cur_gray_reg <= {ADDR_WIDTH+1{1'b0}};

            wr_ptr_update_valid_reg <= 1'b0;
            wr_ptr_update_reg <= 1'b0;
        end
    end
end

// pointer synchronization
always @(posedge s_clk or negedge s_rst_n) begin
    if (!s_rst_n) begin
        rd_ptr_gray_sync1_reg <= {ADDR_WIDTH+1{1'b0}};
        rd_ptr_gray_sync2_reg <= {ADDR_WIDTH+1{1'b0}};
        wr_ptr_update_ack_sync1_reg <= 1'b0;
        wr_ptr_update_ack_sync2_reg <= 1'b0;
    end else begin
        rd_ptr_gray_sync1_reg <= rd_ptr_gray_reg;
        rd_ptr_gray_sync2_reg <= rd_ptr_gray_sync1_reg;
        wr_ptr_update_ack_sync1_reg <= wr_ptr_update_sync3_reg;
        wr_ptr_update_ack_sync2_reg <= wr_ptr_update_ack_sync1_reg;
    end
end

always @(posedge m_clk or negedge m_rst_n) begin
    if (!m_rst_n) begin
        wr_ptr_gray_sync1_reg <= {ADDR_WIDTH+1{1'b0}};
        wr_ptr_gray_sync2_reg <= {ADDR_WIDTH+1{1'b0}};
        wr_ptr_update_sync1_reg <= 1'b0;
        wr_ptr_update_sync2_reg <= 1'b0;
        wr_ptr_update_sync3_reg <= 1'b0;
    end else begin
        if (!FRAME_FIFO) begin
            wr_ptr_gray_sync1_reg <= wr_ptr_gray_reg;
        end else if (wr_ptr_update_sync2_reg ^ wr_ptr_update_sync3_reg) begin
            wr_ptr_gray_sync1_reg <= wr_ptr_sync_gray_reg;
        end
        wr_ptr_gray_sync2_reg <= wr_ptr_gray_sync1_reg;
        wr_ptr_update_sync1_reg <= wr_ptr_update_reg;
        wr_ptr_update_sync2_reg <= wr_ptr_update_sync1_reg;
        wr_ptr_update_sync3_reg <= wr_ptr_update_sync2_reg;

        if (FRAME_FIFO && !m_rst_sync3_reg) begin
            wr_ptr_gray_sync1_reg <= {ADDR_WIDTH+1{1'b0}};
        end
    end
end

// status synchronization
always @(posedge s_clk or negedge s_rst_n) begin
    if (!s_rst_n) begin
        overflow_sync1_reg <= 1'b0;
        bad_frame_sync1_reg <= 1'b0;
        good_frame_sync1_reg <= 1'b0;
    end else begin
        overflow_sync1_reg <= overflow_sync1_reg ^ overflow_reg;
        bad_frame_sync1_reg <= bad_frame_sync1_reg ^ bad_frame_reg;
        good_frame_sync1_reg <= good_frame_sync1_reg ^ good_frame_reg;
    end
end

always @(posedge m_clk or negedge m_rst_n) begin
    if (!m_rst_n) begin
        overflow_sync2_reg <= 1'b0;
        overflow_sync3_reg <= 1'b0;
        overflow_sync4_reg <= 1'b0;
        bad_frame_sync2_reg <= 1'b0;
        bad_frame_sync3_reg <= 1'b0;
        bad_frame_sync4_reg <= 1'b0;
        good_frame_sync2_reg <= 1'b0;
        good_frame_sync3_reg <= 1'b0;
        good_frame_sync4_reg <= 1'b0;
    end else begin
        overflow_sync2_reg <= overflow_sync1_reg;
        overflow_sync3_reg <= overflow_sync2_reg;
        overflow_sync4_reg <= overflow_sync3_reg;
        bad_frame_sync2_reg <= bad_frame_sync1_reg;
        bad_frame_sync3_reg <= bad_frame_sync2_reg;
        bad_frame_sync4_reg <= bad_frame_sync3_reg;
        good_frame_sync2_reg <= good_frame_sync1_reg;
        good_frame_sync3_reg <= good_frame_sync2_reg;
        good_frame_sync4_reg <= good_frame_sync3_reg;
    end
end

// Read logic
integer j;

`ifdef TARGET_XILINX
always @(posedge m_clk) begin // Vivado could not infer BRAM if async reset is used.
`else
always @(posedge m_clk or negedge m_rst_n) begin
`endif
    if (!m_rst_n) begin
        rd_ptr_reg <= {ADDR_WIDTH+1{1'b0}};
        rd_ptr_gray_reg <= {ADDR_WIDTH+1{1'b0}};
        for (j=0; j<PIPELINE_OUTPUT; j=j+1) m_axis_pipe_reg[j] <= 0;
        m_axis_tvalid_pipe_reg <= {PIPELINE_OUTPUT{1'b0}};
        m_frame_reg <= 1'b0;
        m_drop_frame_reg <= 1'b0;
        m_terminate_frame_reg <= 1'b0;
    end else begin
        if (m_axis_tready) begin
            // output ready; invalidate stage
            m_axis_tvalid_pipe_reg[PIPELINE_OUTPUT-1] <= 1'b0;
            m_terminate_frame_reg <= 1'b0;
        end

        for (j = PIPELINE_OUTPUT-1; j > 0; j = j - 1) begin
            if (m_axis_tready || |((~m_axis_tvalid_pipe_reg) >> j)) begin
                // output ready or bubble in pipeline; transfer down pipeline
                m_axis_tvalid_pipe_reg[j] <= m_axis_tvalid_pipe_reg[j-1];
                m_axis_pipe_reg[j] <= m_axis_pipe_reg[j-1];
                m_axis_tvalid_pipe_reg[j-1] <= 1'b0;
            end
        end

        if (m_axis_tready || |(~m_axis_tvalid_pipe_reg)) begin
            // output ready or bubble in pipeline; read new data from FIFO
            m_axis_tvalid_pipe_reg[0] <= 1'b0;
            m_axis_pipe_reg[0] <= mem[rd_ptr_reg[ADDR_WIDTH-1:0]];
            if (!empty && m_rst_sync3_reg && !m_drop_frame_reg) begin
                // not empty, increment pointer
                m_axis_tvalid_pipe_reg[0] <= 1'b1;
                rd_ptr_reg <= rd_ptr_reg + 1;
                rd_ptr_gray_reg <= (rd_ptr_reg + 1) ^ ((rd_ptr_reg + 1) >> 1);
            end
        end

        if (m_axis_tvalid && LAST_ENABLE) begin
            // track output frame status
            if (m_axis_tlast && m_axis_tready) begin
                m_frame_reg <= 1'b0;
            end else begin
                m_frame_reg <= 1'b1;
            end
        end

        if (m_drop_frame_reg && (m_axis_tready || !m_axis_tvalid_pipe) && LAST_ENABLE) begin
            // terminate frame
            // (only for frame transfers interrupted by source reset)
            m_axis_tvalid_pipe_reg[PIPELINE_OUTPUT-1] <= 1'b1;
            m_terminate_frame_reg <= 1'b1;
            m_drop_frame_reg <= 1'b0;
        end

        if (!m_rst_sync3_reg && LAST_ENABLE) begin
            // if source side is reset during transfer, drop partial frame

            // empty output pipeline, except for last stage
            if (PIPELINE_OUTPUT > 1) begin
                m_axis_tvalid_pipe_reg[PIPELINE_OUTPUT-2:0] <= 0;
            end

            if (m_frame_reg && (!m_axis_tvalid || (m_axis_tvalid && !m_axis_tlast)) &&
                    !(m_drop_frame_reg || m_terminate_frame_reg)) begin
                // terminate frame
                m_drop_frame_reg <= 1'b1;
            end
        end

        if (!m_rst_sync3_reg) begin
            rd_ptr_reg <= {ADDR_WIDTH+1{1'b0}};
            rd_ptr_gray_reg <= {ADDR_WIDTH+1{1'b0}};
        end
    end
end

endmodule

`resetall
