`define IP_HDR_SIZE 20
`define
`define IP_HDR_OFFSET_VERSION_IHL 0  // Version, IHL
`define IP_HDR_OFFSET_TOS         1  // Type of Service
`define IP_HDR_OFFSET_TOT_LEN     2  // Total Length
`define IP_HDR_OFFSET_ID          4  // Identification
`define IP_HDR_OFFSET_FLAG_OFF    6  // Flags, Fragment Offset
`define IP_HDR_OFFSET_TTL         8  // Time to Live
`define IP_HDR_OFFSET_PROTOCOL    9  // Protocol
`define IP_HDR_OFFSET_CHECK       10 // Header Checksum
`define IP_HDR_OFFSET_SADDR       12 // Source Address
`define IP_HDR_OFFSET_DADDR       16 // Destination Address
